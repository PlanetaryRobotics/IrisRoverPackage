
module read_register_table(/* from the intr_data_buffer */
							 input [7:0]   reg_addr,
							 input [127:0] reg_data,
							 input         valid_reg_stuff,
							 
							 
							 output 
							 
							 
							 
							
							 
							 