module FPGA_Interpolation_JPG_Block(input sysClk,
												input[11:0] dozen_in,
												input metadata_flag,
												input pixeldata_flag,
												
												output byte_to_store,
												output valid_byte_flag
												);
												
			
endmodule