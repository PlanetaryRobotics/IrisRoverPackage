module bayer_interpolation(input sysClk,
													 input[11:0] bayer_image_in[1943:0][2591:0],
													 input input_valid,

													 output[35:0] RGB_image[1943:0][2591:0],
													 output output_valid);


endmodule
