module bayer_to_rgb(input sysClk,
                    input[11:0]
                    );

endmodule
