module num_img_stored_reg(input[15:0]  in_num_nav_img_numimg_reg,
								  input[31:16] in_num_science_img_numimg_reg,
								  
								  input        in_valid_numimg_reg,
								  
								  input        start_flush_numimg_reg,
								  
								  output[31:0] out_numimg_reg,
								  output		   out_valid_numimg_reg
								  );
								  
								  



endmodule